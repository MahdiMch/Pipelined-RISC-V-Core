`include "Data_mem.v"
module memory_cycle(clk,rst,PCSrcE,RegWriteM,MemWriteM,ResultSrcM,RD_M,PCTargetE,PCPlus4M,WriteDataM,ALU_ResultM,RegWriteW,ResultSrcW,RD_W,PCPlus4W,ALU_ResultW,ReadDataW);
    input clk,rst,PCSrcE,RegWriteM,MemWriteM,ResultSrcM;
    input [4:0] RD_M;
    input [31:0] PCPlus4M,WriteDataM,ALU_ResultM,PCTargetE;
    output RegWriteW,ResultSrcW;
    output [4:0] RD_W;
    output [31:0] PCPlus4W,ALU_ResultW,ReadDataW;

    wire [31:0] ReadDataM;
    reg RegWriteM_r,MemWriteM_r,ResultSrcM_r;
    reg [4:0] RD_M_r;
    reg [31:0] PCPlus4M_r,ReadDataM_r,ALU_ResultM_r;
    Data_mem data_mem(
        .clk(clk),
        .rst(rst),
        .WE(MemWriteM),
        .WD(WriteDataM),
        .A(ALU_ResultM),
        .RD(ReadDataM)
    );
    always @(posedge clk or negedge rst) begin
        if (rst==1'b0) begin
            RegWriteM_r <= 1'b0;
            ResultSrcM_r <= 1'b0;
            RD_M_r <= 5'h00;
            PCPlus4M_r <= 32'h00000000;
            ALU_ResultM_r <= 32'h00000000;
            ReadDataM_r <= 32'h00000000;
        end
        else begin
            RegWriteM_r <= RegWriteM;
            ResultSrcM_r <= MemWriteM;
            RD_M_r <= RD_M;
            PCPlus4M_r <= PCPlus4M;
            ALU_ResultM_r <= ALU_ResultM;
            ReadDataM_r <= ReadDataM;
        end

    end 
assign RegWriteW = RegWriteM_r;
assign ResultSrcW = ResultSrcM_r;
assign RD_W = RD_M_r;
assign PCPlus4W = PCPlus4M_r;
assign ALU_ResultW = ALU_ResultM_r;
assign ReadDataW = ReadDataM_r;


endmodule